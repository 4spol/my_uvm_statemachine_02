interface my_ifo (input  clk,input  rst_n) ;//the dut  output interface
	logic en;
	logic [2:0]cnt;
	logic vaild;
endinterface

