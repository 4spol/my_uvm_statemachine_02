class base_test extends uvm_test;//base_test for other test extending

   my_env         env;
   
   function new(string name = "base_test", uvm_component parent = null);
      super.new(name,parent);
   endfunction
   
   extern virtual function void build_phase(uvm_phase phase);
   extern virtual task  main_phase(uvm_phase phase);
   extern virtual function void report_phase(uvm_phase phase);
   `uvm_component_utils(base_test)
endclass


function void base_test::build_phase(uvm_phase phase);
   super.build_phase(phase);
   env  =  my_env::type_id::create("env", this); //new env
endfunction

task  base_test::main_phase(uvm_phase phase);
   phase.phase_done.set_drain_time(this,200);//set_drain_time for monitoro to get info
endtask

function void base_test::report_phase(uvm_phase phase);//check error number
   uvm_report_server server;
   int err_num;
   super.report_phase(phase);
   server = get_report_server();
   err_num = server.get_severity_count(UVM_ERROR);

   if (err_num != 0) begin
      $display("TEST CASE FAILED");
   end
   else begin
      $display("TEST CASE PASSED");
   end
endfunction


