interface my_if (input  clk,input  rst_n);//the dut input interface
	logic  vaild;
	logic  data;
endinterface


